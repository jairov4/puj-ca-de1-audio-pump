module avl_mm_master_export
(clk, reset,
avm_readdata, avm_writedata, avm_read, avm_write, avm_address, avm_waitrequest,
e_readdata, e_writedata, e_read, e_write, e_address, e_waitrequest, clk, reset);


endmodule;